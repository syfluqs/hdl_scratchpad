-- can_master_coord.vhdl
-- author: roy
-- created: 2017-10-24
-- description : coordinates the can bus masters, acts like a testbench

library ieee;
use ieee.std_logic_1164.all;

